library verilog;
use verilog.vl_types.all;
entity sim_fifo_top is
    generic(
        DATA_WIDTH      : integer := 32;
        DO_WIDTH        : integer := 64;
        BANK_WIDTH      : integer := 3;
        CKE_WIDTH       : integer := 1;
        CLK_WIDTH       : integer := 4;
        COL_WIDTH       : integer := 10;
        CS_NUM          : integer := 1;
        CS_WIDTH        : integer := 4;
        CS_BITS         : integer := 0;
        DQ_WIDTH        : integer := 32;
        DM_WIDTH        : integer := 4;
        DQ_PER_DQS      : integer := 8;
        DQS_WIDTH       : integer := 4;
        DQ_BITS         : integer := 5;
        DQS_BITS        : integer := 2;
        ODT_WIDTH       : integer := 4;
        ROW_WIDTH       : integer := 15;
        ADDITIVE_LAT    : integer := 0;
        BURST_LEN       : integer := 8;
        BURST_TYPE      : integer := 0;
        CAS_LAT         : integer := 4;
        ECC_ENABLE      : integer := 0;
        APPDATA_WIDTH   : integer := 64;
        MULTI_BANK_EN   : integer := 1;
        TWO_T_TIME_EN   : integer := 0;
        ODT_TYPE        : integer := 1;
        REDUCE_DRV      : integer := 0;
        REG_ENABLE      : integer := 0;
        TREFI_NS        : integer := 7800;
        TRAS            : integer := 40000;
        TRCD            : integer := 15000;
        TRFC            : integer := 197500;
        TRP             : integer := 15000;
        TRTP            : integer := 7500;
        TWR             : integer := 15000;
        TWTR            : integer := 7500;
        HIGH_PERFORMANCE_MODE: string  := "TRUE";
        SIM_ONLY        : integer := 0;
        DEBUG_EN        : integer := 0;
        CLK_PERIOD      : integer := 3750;
        DLL_FREQ_MODE   : string  := "HIGH";
        CLK_TYPE        : string  := "SINGLE_ENDED";
        NOCLK200        : integer := 0;
        RST_ACT_LOW     : integer := 1
    );
    port(
        data_in         : in     vl_logic_vector;
        wr_clk          : in     vl_logic;
        ref_clk         : in     vl_logic;
        sys_clk         : in     vl_logic;
        clk_200         : in     vl_logic;
        rd_clk          : in     vl_logic;
        reset_n         : in     vl_logic;
        wr_en           : in     vl_logic;
        rd_en           : in     vl_logic;
        full            : out    vl_logic;
        almost_full     : out    vl_logic;
        empty           : out    vl_logic;
        almost_empty    : out    vl_logic;
        phy_init_done   : out    vl_logic;
        dout_vd         : out    vl_logic;
        data_out        : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DO_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CLK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CS_NUM : constant is 1;
    attribute mti_svvh_generic_type of CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CS_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQ_PER_DQS : constant is 1;
    attribute mti_svvh_generic_type of DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQ_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQS_BITS : constant is 1;
    attribute mti_svvh_generic_type of ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ADDITIVE_LAT : constant is 1;
    attribute mti_svvh_generic_type of BURST_LEN : constant is 1;
    attribute mti_svvh_generic_type of BURST_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CAS_LAT : constant is 1;
    attribute mti_svvh_generic_type of ECC_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of APPDATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MULTI_BANK_EN : constant is 1;
    attribute mti_svvh_generic_type of TWO_T_TIME_EN : constant is 1;
    attribute mti_svvh_generic_type of ODT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of REDUCE_DRV : constant is 1;
    attribute mti_svvh_generic_type of REG_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TREFI_NS : constant is 1;
    attribute mti_svvh_generic_type of TRAS : constant is 1;
    attribute mti_svvh_generic_type of TRCD : constant is 1;
    attribute mti_svvh_generic_type of TRFC : constant is 1;
    attribute mti_svvh_generic_type of TRP : constant is 1;
    attribute mti_svvh_generic_type of TRTP : constant is 1;
    attribute mti_svvh_generic_type of TWR : constant is 1;
    attribute mti_svvh_generic_type of TWTR : constant is 1;
    attribute mti_svvh_generic_type of HIGH_PERFORMANCE_MODE : constant is 1;
    attribute mti_svvh_generic_type of SIM_ONLY : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_EN : constant is 1;
    attribute mti_svvh_generic_type of CLK_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of DLL_FREQ_MODE : constant is 1;
    attribute mti_svvh_generic_type of CLK_TYPE : constant is 1;
    attribute mti_svvh_generic_type of NOCLK200 : constant is 1;
    attribute mti_svvh_generic_type of RST_ACT_LOW : constant is 1;
end sim_fifo_top;
